// This is a generated file. Use and modify at your own risk.
//////////////////////////////////////////////////////////////////////////////// 
// default_nettype of none prevents implicit wire declaration.
`default_nettype none
module axonerve_kvs_rtl_example #(
  parameter integer C_M00_AXI_ADDR_WIDTH = 64  ,
  parameter integer C_M00_AXI_DATA_WIDTH = 512
)
(
  // System Signals
  input  wire                              ap_clk         ,
  input  wire                              ap_rst_n       ,
  // AXI4 master interface m00_axi
  output wire                              m00_axi_awvalid,
  input  wire                              m00_axi_awready,
  output wire [C_M00_AXI_ADDR_WIDTH-1:0]   m00_axi_awaddr ,
  output wire [8-1:0]                      m00_axi_awlen  ,
  output wire                              m00_axi_wvalid ,
  input  wire                              m00_axi_wready ,
  output wire [C_M00_AXI_DATA_WIDTH-1:0]   m00_axi_wdata  ,
  output wire [C_M00_AXI_DATA_WIDTH/8-1:0] m00_axi_wstrb  ,
  output wire                              m00_axi_wlast  ,
  input  wire                              m00_axi_bvalid ,
  output wire                              m00_axi_bready ,
  output wire                              m00_axi_arvalid,
  input  wire                              m00_axi_arready,
  output wire [C_M00_AXI_ADDR_WIDTH-1:0]   m00_axi_araddr ,
  output wire [8-1:0]                      m00_axi_arlen  ,
  input  wire                              m00_axi_rvalid ,
  output wire                              m00_axi_rready ,
  input  wire [C_M00_AXI_DATA_WIDTH-1:0]   m00_axi_rdata  ,
  input  wire                              m00_axi_rlast  ,
  // SDx Control Signals
  input  wire                              ap_start       ,
  output wire                              ap_idle        ,
  output wire                              ap_done        ,
  input  wire [32-1:0]                     data_num       ,
  input  wire [64-1:0]                     axi00_ptr0     
);


timeunit 1ps;
timeprecision 1ps;

///////////////////////////////////////////////////////////////////////////////
// Local Parameters
///////////////////////////////////////////////////////////////////////////////
// Large enough for interesting traffic.
localparam integer  LP_DEFAULT_LENGTH_IN_BYTES = 16384;
localparam integer  LP_NUM_EXAMPLES    = 1;

///////////////////////////////////////////////////////////////////////////////
// Wires and Variables
///////////////////////////////////////////////////////////////////////////////
(* KEEP = "yes" *)
logic                                areset                         = 1'b0;
logic                                ap_start_r                     = 1'b0;
logic                                ap_idle_r                      = 1'b1;
logic                                ap_start_pulse                ;
logic [LP_NUM_EXAMPLES-1:0]          ap_done_i                     ;
logic [LP_NUM_EXAMPLES-1:0]          ap_done_r                      = {LP_NUM_EXAMPLES{1'b0}};
logic [32-1:0]                       ctrl_xfer_size_in_bytes        = LP_DEFAULT_LENGTH_IN_BYTES;
logic [32-1:0]                       ctrl_constant                  = 32'd1;

///////////////////////////////////////////////////////////////////////////////
// Begin RTL
///////////////////////////////////////////////////////////////////////////////

//`define SIMULATION

`ifndef SIMULATION
always @(posedge ap_clk) begin
   ctrl_xfer_size_in_bytes <= data_num;
end
`endif

// Register and invert reset signal.
always @(posedge ap_clk) begin
  areset <= ~ap_rst_n;
end

// create pulse when ap_start transitions to 1
always @(posedge ap_clk) begin
  begin
    ap_start_r <= ap_start;
  end
end

assign ap_start_pulse = ap_start & ~ap_start_r;

// ap_idle is asserted when done is asserted, it is de-asserted when ap_start_pulse
// is asserted
always @(posedge ap_clk) begin
  if (areset) begin
    ap_idle_r <= 1'b1;
  end
  else begin
    ap_idle_r <= ap_done ? 1'b1 :
      ap_start_pulse ? 1'b0 : ap_idle;
  end
end

assign ap_idle = ap_idle_r;

// Done logic
always @(posedge ap_clk) begin
  if (areset) begin
    ap_done_r <= '0;
  end
  else begin
    ap_done_r <= (ap_start_pulse | ap_done) ? '0 : ap_done_r | ap_done_i;
  end
end

assign ap_done = &ap_done_r;

   logic clk_100mhz, clk_200mhz;
   logic reset_100mhz = 1'b1;
   logic [7:0] reset_counter_100mhz = 8'd0;

   always @(posedge clk_100mhz) begin
      if(reset_counter_100mhz < 8'd10) begin
	 reset_counter_100mhz <= reset_counter_100mhz + 1;
	 reset_100mhz <= 1'b1;
      end else begin
	 reset_100mhz <= 1'b0;
      end
   end

   clk_wiz_0 inst_clk_wiz_0
     (
      // Clock out ports
      .clk_out1(clk_100mhz),
      .clk_out2(clk_200mhz),
      // Status and control signals
      .reset(areset),
      .locked(),
      .clk_in1(ap_clk)
      );

   logic                            p00_rd_tvalid;
   logic                            p00_rd_tready;
   logic                            p00_rd_tlast;
   logic [C_M00_AXI_DATA_WIDTH-1:0] p00_rd_tdata;
   logic 			    p00_wr_tvalid;
   logic 			    p00_wr_tready;
   logic [C_M00_AXI_DATA_WIDTH-1:0] p00_wr_tdata;
   
// Vadd example
axonerve_kvs_rtl_example_vadd #(
  .C_M_AXI_ADDR_WIDTH ( C_M00_AXI_ADDR_WIDTH ),
  .C_M_AXI_DATA_WIDTH ( C_M00_AXI_DATA_WIDTH ),
  .C_ADDER_BIT_WIDTH  ( 32                   ),
  .C_XFER_SIZE_WIDTH  ( 32                   )
)
inst_example_vadd_m00_axi (
  .aclk                    ( ap_clk                  ),
  .areset                  ( areset                  ),
  .kernel_clk              ( clk_100mhz              ),
  .kernel_rst              ( reset_100mhz            ),
  .ctrl_addr_offset        ( axi00_ptr0              ),
  .ctrl_xfer_size_in_bytes ( ctrl_xfer_size_in_bytes ),
  .ctrl_constant           ( 32'b1                   ),
  .ap_start                ( ap_start_pulse          ),
  .ap_done                 ( ap_done_i[0]            ),
  .m_axi_awvalid           ( m00_axi_awvalid         ),
  .m_axi_awready           ( m00_axi_awready         ),
  .m_axi_awaddr            ( m00_axi_awaddr          ),
  .m_axi_awlen             ( m00_axi_awlen           ),
  .m_axi_wvalid            ( m00_axi_wvalid          ),
  .m_axi_wready            ( m00_axi_wready          ),
  .m_axi_wdata             ( m00_axi_wdata           ),
  .m_axi_wstrb             ( m00_axi_wstrb           ),
  .m_axi_wlast             ( m00_axi_wlast           ),
  .m_axi_bvalid            ( m00_axi_bvalid          ),
  .m_axi_bready            ( m00_axi_bready          ),
  .m_axi_arvalid           ( m00_axi_arvalid         ),
  .m_axi_arready           ( m00_axi_arready         ),
  .m_axi_araddr            ( m00_axi_araddr          ),
  .m_axi_arlen             ( m00_axi_arlen           ),
  .m_axi_rvalid            ( m00_axi_rvalid          ),
  .m_axi_rready            ( m00_axi_rready          ),
  .m_axi_rdata             ( m00_axi_rdata           ),
  .m_axi_rlast             ( m00_axi_rlast           ),

  .rd_tvalid(p00_rd_tvalid),
  .rd_tready(p00_rd_tready),
  .rd_tlast (p00_rd_tlast),
  .rd_tdata (p00_rd_tdata),
  .wr_tvalid(p00_wr_tvalid),
  .wr_tready(p00_wr_tready),
  .wr_tdata (p00_wr_tdata)
			   
);

user_logic #(
	     .C_M_AXI_DATA_WIDTH(C_M00_AXI_DATA_WIDTH)
	     )
   inst_user_logic (
		    .aclk       (ap_clk),
		    .areset     (areset),
		    .kernel_clk (clk_100mhz),
		    .kernel_rst (reset_100mhz),
		    .kernel_clk_2x (clk_200mhz),
    
		    .p00_rd_tvalid(p00_rd_tvalid),
		    .p00_rd_tready(p00_rd_tready),
		    .p00_rd_tlast (p00_rd_tlast),
		    .p00_rd_tdata (p00_rd_tdata),
		    .p00_wr_tvalid(p00_wr_tvalid),
		    .p00_wr_tready(p00_wr_tready),
		    .p00_wr_tdata (p00_wr_tdata)
    );

endmodule : axonerve_kvs_rtl_example
`default_nettype wire
